module m_axia_mem #(
) (
);

endmodule
