module s_axi_mem #(
) (
);

endmodule
