module m_axi_mem #(
) (
);


endmodule
