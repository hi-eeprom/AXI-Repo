module m_axi_mem #(
  parameter SLAVE_BASE_ADDR = 32'h40000000,
  parameter BURST_LEN = 16,
  parameter ID_WIDTH = 1,
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 32,
  parameter AWUSER_WIDTH = 0,
  parameter ARUSER_WIDTH = 0,
  parameter WUSER_WIDTH = 0,
  parameter RUSER_WIDTH = 0,
  parameter BUSER_WIDTH = 0
) (
  input  logic txn_start,
  output logic txn_done,
  output logic txn_error,
  
  input  logic m_axi_aclk,
  input  logic m_axi_aresetn,
  output logic [ID_WIDTH-1:0] m_axi_awid,
  output logic [ADDR_WIDTH-1:0] m_axi_awaddr,
  output logic [7:0] m_axi_awlen,
  output logic [2:0] m_axi_awsize,
  output logic [1:0] m_axi_awburst,
  output logic m_axi_awlock,
  output logic [3:0] m_axi_awcache,
  output logic [2:0] m_axi_awport,
  output logic [3:0] m_axi_awqos,
  output logic [AWUSER_WIDTH-1:0] m_axi_awuser,
  output logic m_axi_awvalid,
  input  logic m_axi_awready,
  output logic [DATA_WIDTH-1:0] m_axi_wdata,
  output logic [DATA_WIDTH/8-1:0] m_axi_wstrb,
  output logic m_axi_wlast,
  output logic [WUSER_WIDTH-1:0] m_axi_wuser,
  output logic m_axi_wvalid,
  input  logic m_axi_wready,
  input  logic [ID_WIDTH-1:0] m_axi_bid,
  input  logic [1:0] m_axi_bresp,
  input  logic [BUSER_WIDTH-1:0] m_axi_buser,
  input  logic m_axi_wvalid,
  output logic m_axi_wready,
  output logic [ID_WIDTH-1:0] m_axi_arid,
  output logic [ADDR_WIDTH-1:0] m_axi_araddr,
  output logic [7:0] m_axi_arlen,
  output logic [2:0] m_axi_arsize,
  output logic [1:0] m_axi_arburst,
  output logic m_axi_arlock,
  output logic [3:0] m_axi_arcache,
  output logic [2:0] m_axi_arport,
  output logic [3:0] m_axi_arqos,
  output logic [ARUSER_WIDTH-1:0] m_axi_aruser,
  output logic m_axi_arvalid,
  input  logic m_axi_arready,
  input  logic [ID_WIDTH-1:0] m_axi_rid,
  input  logic [DATA_WIDTH-1:0] m_axi_rdata,
  input  logic [1:0] m_axi_rresp,
  input  logic [RUSER_WIDTH-1:0] m_axi_ruser,
  input  logic m_axi_rvalid,
  output logic m_axi_rready
);


endmodule
