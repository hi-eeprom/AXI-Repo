module s_axi_interrupt #(
) (
);


endmodule
